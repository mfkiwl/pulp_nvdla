`ifndef DESIGNWARE_NOEXIST
    `define DESIGNWARE_NOEXIST
`endif