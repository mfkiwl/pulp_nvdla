`ifndef NVTOOLS_SYNC2D_GENERIC_CELL
    `define NVTOOLS_SYNC2D_GENERIC_CELL
`endif